module fifo_v3_25BB5_2766A (
	clk_i,
	rst_ni,
	flush_i,
	testmode_i,
	full_o,
	empty_o,
	usage_o,
	data_i,
	push_i,
	data_o,
	pop_i
);
	parameter [31:0] dtype_T_AddrWidth = 0;
	parameter [31:0] dtype_T_DataWidth = 0;
	parameter [31:0] dtype_T_IdWidth = 0;
	parameter [31:0] dtype_T_UserWidth = 0;
	reg _sv2v_0;
	parameter [0:0] FALL_THROUGH = 1'b0;
	parameter [31:0] DATA_WIDTH = 32;
	parameter [31:0] DEPTH = 8;
	parameter [31:0] ADDR_DEPTH = (DEPTH > 1 ? $clog2(DEPTH) : 1);
	input wire clk_i;
	input wire rst_ni;
	input wire flush_i;
	input wire testmode_i;
	output wire full_o;
	output wire empty_o;
	output wire [ADDR_DEPTH - 1:0] usage_o;
	input wire [(((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10:0] data_i;
	input wire push_i;
	output reg [(((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10:0] data_o;
	input wire pop_i;
	localparam [31:0] FifoDepth = (DEPTH > 0 ? DEPTH : 1);
	reg gate_clock;
	reg [ADDR_DEPTH - 1:0] read_pointer_n;
	reg [ADDR_DEPTH - 1:0] read_pointer_q;
	reg [ADDR_DEPTH - 1:0] write_pointer_n;
	reg [ADDR_DEPTH - 1:0] write_pointer_q;
	reg [ADDR_DEPTH:0] status_cnt_n;
	reg [ADDR_DEPTH:0] status_cnt_q;
	reg [(((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? (FifoDepth * ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 11)) - 1 : (FifoDepth * (1 - ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10))) + ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 9)):(((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? 0 : (((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10)] mem_n;
	reg [(((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? (FifoDepth * ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 11)) - 1 : (FifoDepth * (1 - ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10))) + ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 9)):(((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? 0 : (((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10)] mem_q;
	assign usage_o = status_cnt_q[ADDR_DEPTH - 1:0];
	generate
		if (DEPTH == 0) begin : gen_pass_through
			assign empty_o = ~push_i;
			assign full_o = ~pop_i;
		end
		else begin : gen_fifo
			assign full_o = status_cnt_q == FifoDepth[ADDR_DEPTH:0];
			assign empty_o = (status_cnt_q == 0) & ~(FALL_THROUGH & push_i);
		end
	endgenerate
	always @(*) begin : read_write_comb
		if (_sv2v_0)
			;
		read_pointer_n = read_pointer_q;
		write_pointer_n = write_pointer_q;
		status_cnt_n = status_cnt_q;
		data_o = (DEPTH == 0 ? data_i : mem_q[(((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? 0 : (((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) + (read_pointer_q * (((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? (((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 11 : 1 - ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10)))+:(((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? (((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 11 : 1 - ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10))]);
		mem_n = mem_q;
		gate_clock = 1'b1;
		if (push_i && ~full_o) begin
			mem_n[(((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? 0 : (((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) + (write_pointer_q * (((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? (((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 11 : 1 - ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10)))+:(((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? (((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 11 : 1 - ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10))] = data_i;
			gate_clock = 1'b0;
			if (write_pointer_q == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				write_pointer_n = 1'sb0;
			else
				write_pointer_n = write_pointer_q + 1;
			status_cnt_n = status_cnt_q + 1;
		end
		if (pop_i && ~empty_o) begin
			if (read_pointer_n == (FifoDepth[ADDR_DEPTH - 1:0] - 1))
				read_pointer_n = 1'sb0;
			else
				read_pointer_n = read_pointer_q + 1;
			status_cnt_n = status_cnt_q - 1;
		end
		if (((push_i && pop_i) && ~full_o) && ~empty_o)
			status_cnt_n = status_cnt_q;
		if ((FALL_THROUGH && (status_cnt_q == 0)) && push_i) begin
			data_o = data_i;
			if (pop_i) begin
				status_cnt_n = status_cnt_q;
				read_pointer_n = read_pointer_q;
				write_pointer_n = write_pointer_q;
			end
		end
	end
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else if (flush_i) begin
			read_pointer_q <= 1'sb0;
			write_pointer_q <= 1'sb0;
			status_cnt_q <= 1'sb0;
		end
		else begin
			read_pointer_q <= read_pointer_n;
			write_pointer_q <= write_pointer_n;
			status_cnt_q <= status_cnt_n;
		end
	function automatic [(((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? (((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 11 : 1 - ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10)) - 1:0] sv2v_cast_AEA95;
		input reg [(((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10) >= 0 ? (((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 11 : 1 - ((((((dtype_T_AddrWidth + 7) + (dtype_T_DataWidth / 8)) + dtype_T_IdWidth) + 9) + dtype_T_UserWidth) + 10)) - 1:0] inp;
		sv2v_cast_AEA95 = inp;
	endfunction
	always @(posedge clk_i or negedge rst_ni)
		if (~rst_ni)
			mem_q <= {FifoDepth {sv2v_cast_AEA95(1'sb0)}};
		else if (!gate_clock)
			mem_q <= mem_n;
	initial _sv2v_0 = 0;
endmodule
