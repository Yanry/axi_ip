module axi_fifo_2DE1F_D0182 (
	clk_i,
	rst_ni,
	test_i,
	slv_req_i,
	slv_resp_o,
	mst_req_o,
	mst_resp_i
);
	parameter [31:0] ar_chan_t_IdWidth = 0;
	parameter [31:0] ar_chan_t_MemAddrWidth = 0;
	parameter [31:0] ar_chan_t_UserWidth = 0;
	parameter [31:0] aw_chan_t_IdWidth = 0;
	parameter [31:0] aw_chan_t_MemAddrWidth = 0;
	parameter [31:0] aw_chan_t_UserWidth = 0;
	parameter [31:0] axi_req_t_DataWidth = 0;
	parameter [31:0] axi_req_t_IdWidth = 0;
	parameter [31:0] axi_req_t_MemAddrWidth = 0;
	parameter [31:0] axi_req_t_UserWidth = 0;
	parameter [31:0] axi_resp_t_DataWidth = 0;
	parameter [31:0] axi_resp_t_IdWidth = 0;
	parameter [31:0] axi_resp_t_UserWidth = 0;
	parameter [31:0] b_chan_t_IdWidth = 0;
	parameter [31:0] b_chan_t_UserWidth = 0;
	parameter [31:0] r_chan_t_DataWidth = 0;
	parameter [31:0] r_chan_t_IdWidth = 0;
	parameter [31:0] r_chan_t_UserWidth = 0;
	parameter [31:0] w_chan_t_DataWidth = 0;
	parameter [31:0] w_chan_t_UserWidth = 0;
	parameter [31:0] Depth = 32'd1;
	parameter [0:0] FallThrough = 1'b0;
	input wire clk_i;
	input wire rst_ni;
	input wire test_i;
	input wire [(((((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 35) + axi_req_t_UserWidth) + 1) + (((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth)) + 2) + (((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth)) + 1:0] slv_req_i;
	output wire [(((4 + ((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth)) + 1) + (((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth)) - 1:0] slv_resp_o;
	output wire [(((((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 35) + axi_req_t_UserWidth) + 1) + (((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth)) + 2) + (((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth)) + 1:0] mst_req_o;
	input wire [(((4 + ((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth)) + 1) + (((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth)) - 1:0] mst_resp_i;
	generate
		if (Depth == {32 {1'sb0}}) begin : gen_no_fifo
			assign mst_req_o = slv_req_i;
			assign slv_resp_o = mst_resp_i;
		end
		else begin : gen_axi_fifo
			wire aw_fifo_empty;
			wire ar_fifo_empty;
			wire w_fifo_empty;
			wire r_fifo_empty;
			wire b_fifo_empty;
			wire aw_fifo_full;
			wire ar_fifo_full;
			wire w_fifo_full;
			wire r_fifo_full;
			wire b_fifo_full;
			assign mst_req_o[1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)))] = ~aw_fifo_empty;
			assign mst_req_o[1] = ~ar_fifo_empty;
			assign mst_req_o[2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)] = ~w_fifo_empty;
			assign slv_resp_o[(((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0] = ~r_fifo_empty;
			assign slv_resp_o[1 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))] = ~b_fifo_empty;
			assign slv_resp_o[4 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))] = ~aw_fifo_full;
			assign slv_resp_o[3 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))] = ~ar_fifo_full;
			assign slv_resp_o[2 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))] = ~w_fifo_full;
			assign mst_req_o[0] = ~r_fifo_full;
			assign mst_req_o[1 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)] = ~b_fifo_full;
			fifo_v3_F0013_F5619 #(
				.dtype_aw_chan_t_IdWidth(aw_chan_t_IdWidth),
				.dtype_aw_chan_t_MemAddrWidth(aw_chan_t_MemAddrWidth),
				.dtype_aw_chan_t_UserWidth(aw_chan_t_UserWidth),
				.DEPTH(Depth),
				.FALL_THROUGH(FallThrough)
			) i_aw_fifo(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.testmode_i(test_i),
				.full_o(aw_fifo_full),
				.empty_o(aw_fifo_empty),
				.usage_o(),
				.data_i(slv_req_i[(((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 35) + axi_req_t_UserWidth) + (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))))-:(((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 35) + axi_req_t_UserWidth) + (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))))) >= (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2)))) ? (((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 35) + axi_req_t_UserWidth) + (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))))) - (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2))))) + 1 : ((1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2)))) - ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 35) + axi_req_t_UserWidth) + (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)))))) + 1)]),
				.push_i(slv_req_i[1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)))] && slv_resp_o[4 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))]),
				.data_o(mst_req_o[(((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 35) + axi_req_t_UserWidth) + (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))))-:(((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 35) + axi_req_t_UserWidth) + (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))))) >= (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2)))) ? (((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 35) + axi_req_t_UserWidth) + (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))))) - (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2))))) + 1 : ((1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2)))) - ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 35) + axi_req_t_UserWidth) + (1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)))))) + 1)]),
				.pop_i(mst_req_o[1 + ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)))] && mst_resp_i[4 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))])
			);
			fifo_v3_748B1_E8360 #(
				.dtype_ar_chan_t_IdWidth(ar_chan_t_IdWidth),
				.dtype_ar_chan_t_MemAddrWidth(ar_chan_t_MemAddrWidth),
				.dtype_ar_chan_t_UserWidth(ar_chan_t_UserWidth),
				.DEPTH(Depth),
				.FALL_THROUGH(FallThrough)
			) i_ar_fifo(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.testmode_i(test_i),
				.full_o(ar_fifo_full),
				.empty_o(ar_fifo_empty),
				.usage_o(),
				.data_i(slv_req_i[(((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1-:(((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1) >= 2 ? (((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 0 : 3 - ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))]),
				.push_i(slv_req_i[1] && slv_resp_o[3 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))]),
				.data_o(mst_req_o[(((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1-:(((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1) >= 2 ? (((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 0 : 3 - ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))]),
				.pop_i(mst_req_o[1] && mst_resp_i[3 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))])
			);
			fifo_v3_6EF76_12046 #(
				.dtype_w_chan_t_DataWidth(w_chan_t_DataWidth),
				.dtype_w_chan_t_UserWidth(w_chan_t_UserWidth),
				.DEPTH(Depth),
				.FALL_THROUGH(FallThrough)
			) i_w_fifo(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.testmode_i(test_i),
				.full_o(w_fifo_full),
				.empty_o(w_fifo_empty),
				.usage_o(),
				.data_i(slv_req_i[(((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))-:(((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))) >= (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2)) ? (((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))) - (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2))) + 1 : ((2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2)) - ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)))) + 1)]),
				.push_i(slv_req_i[2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)] && slv_resp_o[2 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))]),
				.data_o(mst_req_o[(((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))-:(((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))) >= (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2)) ? (((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1))) - (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2))) + 1 : ((2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 2)) - ((((axi_req_t_DataWidth + (axi_req_t_DataWidth / 8)) + 1) + axi_req_t_UserWidth) + (2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)))) + 1)]),
				.pop_i(mst_req_o[2 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)] && mst_resp_i[2 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))])
			);
			fifo_v3_5C2E3_C6A7B #(
				.dtype_r_chan_t_DataWidth(r_chan_t_DataWidth),
				.dtype_r_chan_t_IdWidth(r_chan_t_IdWidth),
				.dtype_r_chan_t_UserWidth(r_chan_t_UserWidth),
				.DEPTH(Depth),
				.FALL_THROUGH(FallThrough)
			) i_r_fifo(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.testmode_i(test_i),
				.full_o(r_fifo_full),
				.empty_o(r_fifo_empty),
				.usage_o(),
				.data_i(mst_resp_i[(((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) - 1-:((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth]),
				.push_i(mst_resp_i[(((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0] && mst_req_o[0]),
				.data_o(slv_resp_o[(((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) - 1-:((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth]),
				.pop_i(slv_resp_o[(((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0] && slv_req_i[0])
			);
			fifo_v3_5F756_B22CA #(
				.dtype_b_chan_t_IdWidth(b_chan_t_IdWidth),
				.dtype_b_chan_t_UserWidth(b_chan_t_UserWidth),
				.DEPTH(Depth),
				.FALL_THROUGH(FallThrough)
			) i_b_fifo(
				.clk_i(clk_i),
				.rst_ni(rst_ni),
				.flush_i(1'b0),
				.testmode_i(test_i),
				.full_o(b_fifo_full),
				.empty_o(b_fifo_empty),
				.usage_o(),
				.data_i(mst_resp_i[((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0)-:((((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0)) >= (1 + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0)) ? ((((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0)) - (1 + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))) + 1 : ((1 + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0)) - (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))) + 1)]),
				.push_i(mst_resp_i[1 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))] && mst_req_o[1 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)]),
				.data_o(slv_resp_o[((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0)-:((((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0)) >= (1 + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0)) ? ((((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0)) - (1 + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))) + 1 : ((1 + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0)) - (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))) + 1)]),
				.pop_i(slv_resp_o[1 + (((axi_resp_t_IdWidth + 2) + axi_resp_t_UserWidth) + ((((axi_resp_t_IdWidth + axi_resp_t_DataWidth) + 3) + axi_resp_t_UserWidth) + 0))] && slv_req_i[1 + ((((axi_req_t_IdWidth + axi_req_t_MemAddrWidth) + 29) + axi_req_t_UserWidth) + 1)])
			);
		end
	endgenerate
endmodule
